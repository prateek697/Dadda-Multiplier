`timescale 1ns / 1ps


module adder64bit
(
  input [63:0] x,
  input [63:0] y,
  output [63:0] s
);

 
  wire c0, c1, c2, c3, c4, c5, c6, c7, c8, c9, c10;
  wire c11, c12, c13, c14, c15, c16, c17, c18, c19, c20;
  wire c21, c22, c23, c24, c25, c26, c27, c28, c29, c30;
  wire c31, c32, c33, c34, c35, c36, c37, c38, c39, c40;
  wire c41, c42, c43, c44, c45, c46, c47, c48, c49, c50;
  wire c51, c52, c53, c54, c55, c56, c57, c58, c59, c60;
  wire c61, c62, c63;

 
  assign c0 = 1'b0;

 
  FA k1 (x[0], y[0], c0, s[0], c1);
  FA k2 (x[1], y[1], c1, s[1], c2);
  FA k3 (x[2], y[2], c2, s[2], c3);
  FA k4 (x[3], y[3], c3, s[3], c4);
  FA k5 (x[4], y[4], c4, s[4], c5);
  FA k6 (x[5], y[5], c5, s[5], c6);
  FA k7 (x[6], y[6], c6, s[6], c7);
  FA k8 (x[7], y[7], c7, s[7], c8);
  FA k9 (x[8], y[8], c8, s[8], c9);
  FA k10 (x[9], y[9], c9, s[9], c10);
  FA k11 (x[10], y[10], c10, s[10], c11);
  FA k12 (x[11], y[11], c11, s[11], c12);
  FA k13 (x[12], y[12], c12, s[12], c13);
  FA k14 (x[13], y[13], c13, s[13], c14);
  FA k15 (x[14], y[14], c14, s[14], c15);
  FA k16 (x[15], y[15], c15, s[15], c16);
  FA k17 (x[16], y[16], c16, s[16], c17);
  FA k18 (x[17], y[17], c17, s[17], c18);
  FA k19 (x[18], y[18], c18, s[18], c19);
  FA k20 (x[19], y[19], c19, s[19], c20);
  FA k21 (x[20], y[20], c20, s[20], c21);
  FA k22 (x[21], y[21], c21, s[21], c22);
  FA k23 (x[22], y[22], c22, s[22], c23);
  FA k24 (x[23], y[23], c23, s[23], c24);
  FA k25 (x[24], y[24], c24, s[24], c25);
  FA k26 (x[25], y[25], c25, s[25], c26);
  FA k27 (x[26], y[26], c26, s[26], c27);
  FA k28 (x[27], y[27], c27, s[27], c28);
  FA k29 (x[28], y[28], c28, s[28], c29);
  FA k30 (x[29], y[29], c29, s[29], c30);
  FA k31 (x[30], y[30], c30, s[30], c31);
  FA k32 (x[31], y[31], c31, s[31], c32);
  FA k33 (x[32], y[32], c32, s[32], c33);
  FA k34 (x[33], y[33], c33, s[33], c34);
  FA k35 (x[34], y[34], c34, s[34], c35);
  FA k36 (x[35], y[35], c35, s[35], c36);
  FA k37 (x[36], y[36], c36, s[36], c37);
  FA k38 (x[37], y[37], c37, s[37], c38);
  FA k39 (x[38], y[38], c38, s[38], c39);
  FA k40 (x[39], y[39], c39, s[39], c40);
  FA k41 (x[40], y[40], c40, s[40], c41);
  FA k42 (x[41], y[41], c41, s[41], c42);
  FA k43 (x[42], y[42], c42, s[42], c43);
  FA k44 (x[43], y[43], c43, s[43], c44);
  FA k45 (x[44], y[44], c44, s[44], c45);
  FA k46 (x[45], y[45], c45, s[45], c46);
  FA k47 (x[46], y[46], c46, s[46], c47);
  FA k48 (x[47], y[47], c47, s[47], c48);
  FA k49 (x[48], y[48], c48, s[48], c49);
  FA k50 (x[49], y[49], c49, s[49], c50);
  FA k51 (x[50], y[50], c50, s[50], c51);
  FA k52 (x[51], y[51], c51, s[51], c52);
  FA k53 (x[52], y[52], c52, s[52], c53);
  FA k54 (x[53], y[53], c53, s[53], c54);
  FA k55 (x[54], y[54], c54, s[54], c55);
  FA k56 (x[55], y[55], c55, s[55], c56);
  FA k57 (x[56], y[56], c56, s[56], c57);
  FA k58 (x[57], y[57], c57, s[57], c58);
  FA k59 (x[58], y[58], c58, s[58], c59);
  FA k60 (x[59], y[59], c59, s[59], c60);
  FA k61 (x[60], y[60], c60, s[60], c61);
  FA k62 (x[61], y[61], c61, s[61], c62);
  FA k63 (x[62], y[62], c62, s[62], c63);
  FA k64 (x[63], y[63], c63, s[63], c);
endmodule


module FA
(
  input A,
  input B,
  input CARRY_IN,
  output SUM,
  output CARRY_OUT
);

  
  wire tmpSum;
  wire tmp1;
  wire tmp1n;
  wire tmp2;
  wire tmp2n;
  wire tmp3;
  wire tmp4;
  wire tmp5;
  wire tmp6;

  
  xor A1 (tmpSum, A, B);
  xor A2 (SUM, CARRY_IN, tmpSum);

  
  not B1N (tmp1n, B);
  and B1 (tmp1, A, tmp1n);
  not B2N (tmp2n, A);
  and B2 (tmp2, tmp2n, B);
  and B3 (tmp3, A, B);
  and B4 (tmp4, tmp1, CARRY_IN);
  and B5 (tmp5, tmp2, CARRY_IN);
  or B6 (tmp6, tmp4, tmp5);
  or B7 (CARRY_OUT, tmp6, tmp3);
endmodule
module Mult_Wallace32  
(
	input [31:0] x,
	input [31:0] y,
	output [63:0] z
);
assign x = 32'b1010101111111;
assign y = 32'b1010101111111;
wire [31:0] P[31:0];

assign P[0][0] = x[0] & y[0];
assign P[0][1] = x[0] & y[1];
assign P[0][2] = x[0] & y[2];
assign P[0][3] = x[0] & y[3];
assign P[0][4] = x[0] & y[4];
assign P[0][5] = x[0] & y[5];
assign P[0][6] = x[0] & y[6];
assign P[0][7] = x[0] & y[7];
assign P[0][8] = x[0] & y[8];
assign P[0][9] = x[0] & y[9];
assign P[0][10] = x[0] & y[10];
assign P[0][11] = x[0] & y[11];
assign P[0][12] = x[0] & y[12];
assign P[0][13] = x[0] & y[13];
assign P[0][14] = x[0] & y[14];
assign P[0][15] = x[0] & y[15];
assign P[0][16] = x[0] & y[16];
assign P[0][17] = x[0] & y[17];
assign P[0][18] = x[0] & y[18];
assign P[0][19] = x[0] & y[19];
assign P[0][20] = x[0] & y[20];
assign P[0][21] = x[0] & y[21];
assign P[0][22] = x[0] & y[22];
assign P[0][23] = x[0] & y[23];
assign P[0][24] = x[0] & y[24];
assign P[0][25] = x[0] & y[25];
assign P[0][26] = x[0] & y[26];
assign P[0][27] = x[0] & y[27];
assign P[0][28] = x[0] & y[28];
assign P[0][29] = x[0] & y[29];
assign P[0][30] = x[0] & y[30];
assign P[0][31] = x[0] & y[31];
assign P[1][0] = x[1] & y[0];
assign P[1][1] = x[1] & y[1];
assign P[1][2] = x[1] & y[2];
assign P[1][3] = x[1] & y[3];
assign P[1][4] = x[1] & y[4];
assign P[1][5] = x[1] & y[5];
assign P[1][6] = x[1] & y[6];
assign P[1][7] = x[1] & y[7];
assign P[1][8] = x[1] & y[8];
assign P[1][9] = x[1] & y[9];
assign P[1][10] = x[1] & y[10];
assign P[1][11] = x[1] & y[11];
assign P[1][12] = x[1] & y[12];
assign P[1][13] = x[1] & y[13];
assign P[1][14] = x[1] & y[14];
assign P[1][15] = x[1] & y[15];
assign P[1][16] = x[1] & y[16];
assign P[1][17] = x[1] & y[17];
assign P[1][18] = x[1] & y[18];
assign P[1][19] = x[1] & y[19];
assign P[1][20] = x[1] & y[20];
assign P[1][21] = x[1] & y[21];
assign P[1][22] = x[1] & y[22];
assign P[1][23] = x[1] & y[23];
assign P[1][24] = x[1] & y[24];
assign P[1][25] = x[1] & y[25];
assign P[1][26] = x[1] & y[26];
assign P[1][27] = x[1] & y[27];
assign P[1][28] = x[1] & y[28];
assign P[1][29] = x[1] & y[29];
assign P[1][30] = x[1] & y[30];
assign P[1][31] = x[1] & y[31];
assign P[2][0] = x[2] & y[0];
assign P[2][1] = x[2] & y[1];
assign P[2][2] = x[2] & y[2];
assign P[2][3] = x[2] & y[3];
assign P[2][4] = x[2] & y[4];
assign P[2][5] = x[2] & y[5];
assign P[2][6] = x[2] & y[6];
assign P[2][7] = x[2] & y[7];
assign P[2][8] = x[2] & y[8];
assign P[2][9] = x[2] & y[9];
assign P[2][10] = x[2] & y[10];
assign P[2][11] = x[2] & y[11];
assign P[2][12] = x[2] & y[12];
assign P[2][13] = x[2] & y[13];
assign P[2][14] = x[2] & y[14];
assign P[2][15] = x[2] & y[15];
assign P[2][16] = x[2] & y[16];
assign P[2][17] = x[2] & y[17];
assign P[2][18] = x[2] & y[18];
assign P[2][19] = x[2] & y[19];
assign P[2][20] = x[2] & y[20];
assign P[2][21] = x[2] & y[21];
assign P[2][22] = x[2] & y[22];
assign P[2][23] = x[2] & y[23];
assign P[2][24] = x[2] & y[24];
assign P[2][25] = x[2] & y[25];
assign P[2][26] = x[2] & y[26];
assign P[2][27] = x[2] & y[27];
assign P[2][28] = x[2] & y[28];
assign P[2][29] = x[2] & y[29];
assign P[2][30] = x[2] & y[30];
assign P[2][31] = x[2] & y[31];
assign P[3][0] = x[3] & y[0];
assign P[3][1] = x[3] & y[1];
assign P[3][2] = x[3] & y[2];
assign P[3][3] = x[3] & y[3];
assign P[3][4] = x[3] & y[4];
assign P[3][5] = x[3] & y[5];
assign P[3][6] = x[3] & y[6];
assign P[3][7] = x[3] & y[7];
assign P[3][8] = x[3] & y[8];
assign P[3][9] = x[3] & y[9];
assign P[3][10] = x[3] & y[10];
assign P[3][11] = x[3] & y[11];
assign P[3][12] = x[3] & y[12];
assign P[3][13] = x[3] & y[13];
assign P[3][14] = x[3] & y[14];
assign P[3][15] = x[3] & y[15];
assign P[3][16] = x[3] & y[16];
assign P[3][17] = x[3] & y[17];
assign P[3][18] = x[3] & y[18];
assign P[3][19] = x[3] & y[19];
assign P[3][20] = x[3] & y[20];
assign P[3][21] = x[3] & y[21];
assign P[3][22] = x[3] & y[22];
assign P[3][23] = x[3] & y[23];
assign P[3][24] = x[3] & y[24];
assign P[3][25] = x[3] & y[25];
assign P[3][26] = x[3] & y[26];
assign P[3][27] = x[3] & y[27];
assign P[3][28] = x[3] & y[28];
assign P[3][29] = x[3] & y[29];
assign P[3][30] = x[3] & y[30];
assign P[3][31] = x[3] & y[31];
assign P[4][0] = x[4] & y[0];
assign P[4][1] = x[4] & y[1];
assign P[4][2] = x[4] & y[2];
assign P[4][3] = x[4] & y[3];
assign P[4][4] = x[4] & y[4];
assign P[4][5] = x[4] & y[5];
assign P[4][6] = x[4] & y[6];
assign P[4][7] = x[4] & y[7];
assign P[4][8] = x[4] & y[8];
assign P[4][9] = x[4] & y[9];
assign P[4][10] = x[4] & y[10];
assign P[4][11] = x[4] & y[11];
assign P[4][12] = x[4] & y[12];
assign P[4][13] = x[4] & y[13];
assign P[4][14] = x[4] & y[14];
assign P[4][15] = x[4] & y[15];
assign P[4][16] = x[4] & y[16];
assign P[4][17] = x[4] & y[17];
assign P[4][18] = x[4] & y[18];
assign P[4][19] = x[4] & y[19];
assign P[4][20] = x[4] & y[20];
assign P[4][21] = x[4] & y[21];
assign P[4][22] = x[4] & y[22];
assign P[4][23] = x[4] & y[23];
assign P[4][24] = x[4] & y[24];
assign P[4][25] = x[4] & y[25];
assign P[4][26] = x[4] & y[26];
assign P[4][27] = x[4] & y[27];
assign P[4][28] = x[4] & y[28];
assign P[4][29] = x[4] & y[29];
assign P[4][30] = x[4] & y[30];
assign P[4][31] = x[4] & y[31];
assign P[5][0] = x[5] & y[0];
assign P[5][1] = x[5] & y[1];
assign P[5][2] = x[5] & y[2];
assign P[5][3] = x[5] & y[3];
assign P[5][4] = x[5] & y[4];
assign P[5][5] = x[5] & y[5];
assign P[5][6] = x[5] & y[6];
assign P[5][7] = x[5] & y[7];
assign P[5][8] = x[5] & y[8];
assign P[5][9] = x[5] & y[9];
assign P[5][10] = x[5] & y[10];
assign P[5][11] = x[5] & y[11];
assign P[5][12] = x[5] & y[12];
assign P[5][13] = x[5] & y[13];
assign P[5][14] = x[5] & y[14];
assign P[5][15] = x[5] & y[15];
assign P[5][16] = x[5] & y[16];
assign P[5][17] = x[5] & y[17];
assign P[5][18] = x[5] & y[18];
assign P[5][19] = x[5] & y[19];
assign P[5][20] = x[5] & y[20];
assign P[5][21] = x[5] & y[21];
assign P[5][22] = x[5] & y[22];
assign P[5][23] = x[5] & y[23];
assign P[5][24] = x[5] & y[24];
assign P[5][25] = x[5] & y[25];
assign P[5][26] = x[5] & y[26];
assign P[5][27] = x[5] & y[27];
assign P[5][28] = x[5] & y[28];
assign P[5][29] = x[5] & y[29];
assign P[5][30] = x[5] & y[30];
assign P[5][31] = x[5] & y[31];
assign P[6][0] = x[6] & y[0];
assign P[6][1] = x[6] & y[1];
assign P[6][2] = x[6] & y[2];
assign P[6][3] = x[6] & y[3];
assign P[6][4] = x[6] & y[4];
assign P[6][5] = x[6] & y[5];
assign P[6][6] = x[6] & y[6];
assign P[6][7] = x[6] & y[7];
assign P[6][8] = x[6] & y[8];
assign P[6][9] = x[6] & y[9];
assign P[6][10] = x[6] & y[10];
assign P[6][11] = x[6] & y[11];
assign P[6][12] = x[6] & y[12];
assign P[6][13] = x[6] & y[13];
assign P[6][14] = x[6] & y[14];
assign P[6][15] = x[6] & y[15];
assign P[6][16] = x[6] & y[16];
assign P[6][17] = x[6] & y[17];
assign P[6][18] = x[6] & y[18];
assign P[6][19] = x[6] & y[19];
assign P[6][20] = x[6] & y[20];
assign P[6][21] = x[6] & y[21];
assign P[6][22] = x[6] & y[22];
assign P[6][23] = x[6] & y[23];
assign P[6][24] = x[6] & y[24];
assign P[6][25] = x[6] & y[25];
assign P[6][26] = x[6] & y[26];
assign P[6][27] = x[6] & y[27];
assign P[6][28] = x[6] & y[28];
assign P[6][29] = x[6] & y[29];
assign P[6][30] = x[6] & y[30];
assign P[6][31] = x[6] & y[31];
assign P[7][0] = x[7] & y[0];
assign P[7][1] = x[7] & y[1];
assign P[7][2] = x[7] & y[2];
assign P[7][3] = x[7] & y[3];
assign P[7][4] = x[7] & y[4];
assign P[7][5] = x[7] & y[5];
assign P[7][6] = x[7] & y[6];
assign P[7][7] = x[7] & y[7];
assign P[7][8] = x[7] & y[8];
assign P[7][9] = x[7] & y[9];
assign P[7][10] = x[7] & y[10];
assign P[7][11] = x[7] & y[11];
assign P[7][12] = x[7] & y[12];
assign P[7][13] = x[7] & y[13];
assign P[7][14] = x[7] & y[14];
assign P[7][15] = x[7] & y[15];
assign P[7][16] = x[7] & y[16];
assign P[7][17] = x[7] & y[17];
assign P[7][18] = x[7] & y[18];
assign P[7][19] = x[7] & y[19];
assign P[7][20] = x[7] & y[20];
assign P[7][21] = x[7] & y[21];
assign P[7][22] = x[7] & y[22];
assign P[7][23] = x[7] & y[23];
assign P[7][24] = x[7] & y[24];
assign P[7][25] = x[7] & y[25];
assign P[7][26] = x[7] & y[26];
assign P[7][27] = x[7] & y[27];
assign P[7][28] = x[7] & y[28];
assign P[7][29] = x[7] & y[29];
assign P[7][30] = x[7] & y[30];
assign P[7][31] = x[7] & y[31];
assign P[8][0] = x[8] & y[0];
assign P[8][1] = x[8] & y[1];
assign P[8][2] = x[8] & y[2];
assign P[8][3] = x[8] & y[3];
assign P[8][4] = x[8] & y[4];
assign P[8][5] = x[8] & y[5];
assign P[8][6] = x[8] & y[6];
assign P[8][7] = x[8] & y[7];
assign P[8][8] = x[8] & y[8];
assign P[8][9] = x[8] & y[9];
assign P[8][10] = x[8] & y[10];
assign P[8][11] = x[8] & y[11];
assign P[8][12] = x[8] & y[12];
assign P[8][13] = x[8] & y[13];
assign P[8][14] = x[8] & y[14];
assign P[8][15] = x[8] & y[15];
assign P[8][16] = x[8] & y[16];
assign P[8][17] = x[8] & y[17];
assign P[8][18] = x[8] & y[18];
assign P[8][19] = x[8] & y[19];
assign P[8][20] = x[8] & y[20];
assign P[8][21] = x[8] & y[21];
assign P[8][22] = x[8] & y[22];
assign P[8][23] = x[8] & y[23];
assign P[8][24] = x[8] & y[24];
assign P[8][25] = x[8] & y[25];
assign P[8][26] = x[8] & y[26];
assign P[8][27] = x[8] & y[27];
assign P[8][28] = x[8] & y[28];
assign P[8][29] = x[8] & y[29];
assign P[8][30] = x[8] & y[30];
assign P[8][31] = x[8] & y[31];
assign P[9][0] = x[9] & y[0];
assign P[9][1] = x[9] & y[1];
assign P[9][2] = x[9] & y[2];
assign P[9][3] = x[9] & y[3];
assign P[9][4] = x[9] & y[4];
assign P[9][5] = x[9] & y[5];
assign P[9][6] = x[9] & y[6];
assign P[9][7] = x[9] & y[7];
assign P[9][8] = x[9] & y[8];
assign P[9][9] = x[9] & y[9];
assign P[9][10] = x[9] & y[10];
assign P[9][11] = x[9] & y[11];
assign P[9][12] = x[9] & y[12];
assign P[9][13] = x[9] & y[13];
assign P[9][14] = x[9] & y[14];
assign P[9][15] = x[9] & y[15];
assign P[9][16] = x[9] & y[16];
assign P[9][17] = x[9] & y[17];
assign P[9][18] = x[9] & y[18];
assign P[9][19] = x[9] & y[19];
assign P[9][20] = x[9] & y[20];
assign P[9][21] = x[9] & y[21];
assign P[9][22] = x[9] & y[22];
assign P[9][23] = x[9] & y[23];
assign P[9][24] = x[9] & y[24];
assign P[9][25] = x[9] & y[25];
assign P[9][26] = x[9] & y[26];
assign P[9][27] = x[9] & y[27];
assign P[9][28] = x[9] & y[28];
assign P[9][29] = x[9] & y[29];
assign P[9][30] = x[9] & y[30];
assign P[9][31] = x[9] & y[31];
assign P[10][0] = x[10] & y[0];
assign P[10][1] = x[10] & y[1];
assign P[10][2] = x[10] & y[2];
assign P[10][3] = x[10] & y[3];
assign P[10][4] = x[10] & y[4];
assign P[10][5] = x[10] & y[5];
assign P[10][6] = x[10] & y[6];
assign P[10][7] = x[10] & y[7];
assign P[10][8] = x[10] & y[8];
assign P[10][9] = x[10] & y[9];
assign P[10][10] = x[10] & y[10];
assign P[10][11] = x[10] & y[11];
assign P[10][12] = x[10] & y[12];
assign P[10][13] = x[10] & y[13];
assign P[10][14] = x[10] & y[14];
assign P[10][15] = x[10] & y[15];
assign P[10][16] = x[10] & y[16];
assign P[10][17] = x[10] & y[17];
assign P[10][18] = x[10] & y[18];
assign P[10][19] = x[10] & y[19];
assign P[10][20] = x[10] & y[20];
assign P[10][21] = x[10] & y[21];
assign P[10][22] = x[10] & y[22];
assign P[10][23] = x[10] & y[23];
assign P[10][24] = x[10] & y[24];
assign P[10][25] = x[10] & y[25];
assign P[10][26] = x[10] & y[26];
assign P[10][27] = x[10] & y[27];
assign P[10][28] = x[10] & y[28];
assign P[10][29] = x[10] & y[29];
assign P[10][30] = x[10] & y[30];
assign P[10][31] = x[10] & y[31];
assign P[11][0] = x[11] & y[0];
assign P[11][1] = x[11] & y[1];
assign P[11][2] = x[11] & y[2];
assign P[11][3] = x[11] & y[3];
assign P[11][4] = x[11] & y[4];
assign P[11][5] = x[11] & y[5];
assign P[11][6] = x[11] & y[6];
assign P[11][7] = x[11] & y[7];
assign P[11][8] = x[11] & y[8];
assign P[11][9] = x[11] & y[9];
assign P[11][10] = x[11] & y[10];
assign P[11][11] = x[11] & y[11];
assign P[11][12] = x[11] & y[12];
assign P[11][13] = x[11] & y[13];
assign P[11][14] = x[11] & y[14];
assign P[11][15] = x[11] & y[15];
assign P[11][16] = x[11] & y[16];
assign P[11][17] = x[11] & y[17];
assign P[11][18] = x[11] & y[18];
assign P[11][19] = x[11] & y[19];
assign P[11][20] = x[11] & y[20];
assign P[11][21] = x[11] & y[21];
assign P[11][22] = x[11] & y[22];
assign P[11][23] = x[11] & y[23];
assign P[11][24] = x[11] & y[24];
assign P[11][25] = x[11] & y[25];
assign P[11][26] = x[11] & y[26];
assign P[11][27] = x[11] & y[27];
assign P[11][28] = x[11] & y[28];
assign P[11][29] = x[11] & y[29];
assign P[11][30] = x[11] & y[30];
assign P[11][31] = x[11] & y[31];
assign P[12][0] = x[12] & y[0];
assign P[12][1] = x[12] & y[1];
assign P[12][2] = x[12] & y[2];
assign P[12][3] = x[12] & y[3];
assign P[12][4] = x[12] & y[4];
assign P[12][5] = x[12] & y[5];
assign P[12][6] = x[12] & y[6];
assign P[12][7] = x[12] & y[7];
assign P[12][8] = x[12] & y[8];
assign P[12][9] = x[12] & y[9];
assign P[12][10] = x[12] & y[10];
assign P[12][11] = x[12] & y[11];
assign P[12][12] = x[12] & y[12];
assign P[12][13] = x[12] & y[13];
assign P[12][14] = x[12] & y[14];
assign P[12][15] = x[12] & y[15];
assign P[12][16] = x[12] & y[16];
assign P[12][17] = x[12] & y[17];
assign P[12][18] = x[12] & y[18];
assign P[12][19] = x[12] & y[19];
assign P[12][20] = x[12] & y[20];
assign P[12][21] = x[12] & y[21];
assign P[12][22] = x[12] & y[22];
assign P[12][23] = x[12] & y[23];
assign P[12][24] = x[12] & y[24];
assign P[12][25] = x[12] & y[25];
assign P[12][26] = x[12] & y[26];
assign P[12][27] = x[12] & y[27];
assign P[12][28] = x[12] & y[28];
assign P[12][29] = x[12] & y[29];
assign P[12][30] = x[12] & y[30];
assign P[12][31] = x[12] & y[31];
assign P[13][0] = x[13] & y[0];
assign P[13][1] = x[13] & y[1];
assign P[13][2] = x[13] & y[2];
assign P[13][3] = x[13] & y[3];
assign P[13][4] = x[13] & y[4];
assign P[13][5] = x[13] & y[5];
assign P[13][6] = x[13] & y[6];
assign P[13][7] = x[13] & y[7];
assign P[13][8] = x[13] & y[8];
assign P[13][9] = x[13] & y[9];
assign P[13][10] = x[13] & y[10];
assign P[13][11] = x[13] & y[11];
assign P[13][12] = x[13] & y[12];
assign P[13][13] = x[13] & y[13];
assign P[13][14] = x[13] & y[14];
assign P[13][15] = x[13] & y[15];
assign P[13][16] = x[13] & y[16];
assign P[13][17] = x[13] & y[17];
assign P[13][18] = x[13] & y[18];
assign P[13][19] = x[13] & y[19];
assign P[13][20] = x[13] & y[20];
assign P[13][21] = x[13] & y[21];
assign P[13][22] = x[13] & y[22];
assign P[13][23] = x[13] & y[23];
assign P[13][24] = x[13] & y[24];
assign P[13][25] = x[13] & y[25];
assign P[13][26] = x[13] & y[26];
assign P[13][27] = x[13] & y[27];
assign P[13][28] = x[13] & y[28];
assign P[13][29] = x[13] & y[29];
assign P[13][30] = x[13] & y[30];
assign P[13][31] = x[13] & y[31];
assign P[14][0] = x[14] & y[0];
assign P[14][1] = x[14] & y[1];
assign P[14][2] = x[14] & y[2];
assign P[14][3] = x[14] & y[3];
assign P[14][4] = x[14] & y[4];
assign P[14][5] = x[14] & y[5];
assign P[14][6] = x[14] & y[6];
assign P[14][7] = x[14] & y[7];
assign P[14][8] = x[14] & y[8];
assign P[14][9] = x[14] & y[9];
assign P[14][10] = x[14] & y[10];
assign P[14][11] = x[14] & y[11];
assign P[14][12] = x[14] & y[12];
assign P[14][13] = x[14] & y[13];
assign P[14][14] = x[14] & y[14];
assign P[14][15] = x[14] & y[15];
assign P[14][16] = x[14] & y[16];
assign P[14][17] = x[14] & y[17];
assign P[14][18] = x[14] & y[18];
assign P[14][19] = x[14] & y[19];
assign P[14][20] = x[14] & y[20];
assign P[14][21] = x[14] & y[21];
assign P[14][22] = x[14] & y[22];
assign P[14][23] = x[14] & y[23];
assign P[14][24] = x[14] & y[24];
assign P[14][25] = x[14] & y[25];
assign P[14][26] = x[14] & y[26];
assign P[14][27] = x[14] & y[27];
assign P[14][28] = x[14] & y[28];
assign P[14][29] = x[14] & y[29];
assign P[14][30] = x[14] & y[30];
assign P[14][31] = x[14] & y[31];
assign P[15][0] = x[15] & y[0];
assign P[15][1] = x[15] & y[1];
assign P[15][2] = x[15] & y[2];
assign P[15][3] = x[15] & y[3];
assign P[15][4] = x[15] & y[4];
assign P[15][5] = x[15] & y[5];
assign P[15][6] = x[15] & y[6];
assign P[15][7] = x[15] & y[7];
assign P[15][8] = x[15] & y[8];
assign P[15][9] = x[15] & y[9];
assign P[15][10] = x[15] & y[10];
assign P[15][11] = x[15] & y[11];
assign P[15][12] = x[15] & y[12];
assign P[15][13] = x[15] & y[13];
assign P[15][14] = x[15] & y[14];
assign P[15][15] = x[15] & y[15];
assign P[15][16] = x[15] & y[16];
assign P[15][17] = x[15] & y[17];
assign P[15][18] = x[15] & y[18];
assign P[15][19] = x[15] & y[19];
assign P[15][20] = x[15] & y[20];
assign P[15][21] = x[15] & y[21];
assign P[15][22] = x[15] & y[22];
assign P[15][23] = x[15] & y[23];
assign P[15][24] = x[15] & y[24];
assign P[15][25] = x[15] & y[25];
assign P[15][26] = x[15] & y[26];
assign P[15][27] = x[15] & y[27];
assign P[15][28] = x[15] & y[28];
assign P[15][29] = x[15] & y[29];
assign P[15][30] = x[15] & y[30];
assign P[15][31] = x[15] & y[31];
assign P[16][0] = x[16] & y[0];
assign P[16][1] = x[16] & y[1];
assign P[16][2] = x[16] & y[2];
assign P[16][3] = x[16] & y[3];
assign P[16][4] = x[16] & y[4];
assign P[16][5] = x[16] & y[5];
assign P[16][6] = x[16] & y[6];
assign P[16][7] = x[16] & y[7];
assign P[16][8] = x[16] & y[8];
assign P[16][9] = x[16] & y[9];
assign P[16][10] = x[16] & y[10];
assign P[16][11] = x[16] & y[11];
assign P[16][12] = x[16] & y[12];
assign P[16][13] = x[16] & y[13];
assign P[16][14] = x[16] & y[14];
assign P[16][15] = x[16] & y[15];
assign P[16][16] = x[16] & y[16];
assign P[16][17] = x[16] & y[17];
assign P[16][18] = x[16] & y[18];
assign P[16][19] = x[16] & y[19];
assign P[16][20] = x[16] & y[20];
assign P[16][21] = x[16] & y[21];
assign P[16][22] = x[16] & y[22];
assign P[16][23] = x[16] & y[23];
assign P[16][24] = x[16] & y[24];
assign P[16][25] = x[16] & y[25];
assign P[16][26] = x[16] & y[26];
assign P[16][27] = x[16] & y[27];
assign P[16][28] = x[16] & y[28];
assign P[16][29] = x[16] & y[29];
assign P[16][30] = x[16] & y[30];
assign P[16][31] = x[16] & y[31];
assign P[17][0] = x[17] & y[0];
assign P[17][1] = x[17] & y[1];
assign P[17][2] = x[17] & y[2];
assign P[17][3] = x[17] & y[3];
assign P[17][4] = x[17] & y[4];
assign P[17][5] = x[17] & y[5];
assign P[17][6] = x[17] & y[6];
assign P[17][7] = x[17] & y[7];
assign P[17][8] = x[17] & y[8];
assign P[17][9] = x[17] & y[9];
assign P[17][10] = x[17] & y[10];
assign P[17][11] = x[17] & y[11];
assign P[17][12] = x[17] & y[12];
assign P[17][13] = x[17] & y[13];
assign P[17][14] = x[17] & y[14];
assign P[17][15] = x[17] & y[15];
assign P[17][16] = x[17] & y[16];
assign P[17][17] = x[17] & y[17];
assign P[17][18] = x[17] & y[18];
assign P[17][19] = x[17] & y[19];
assign P[17][20] = x[17] & y[20];
assign P[17][21] = x[17] & y[21];
assign P[17][22] = x[17] & y[22];
assign P[17][23] = x[17] & y[23];
assign P[17][24] = x[17] & y[24];
assign P[17][25] = x[17] & y[25];
assign P[17][26] = x[17] & y[26];
assign P[17][27] = x[17] & y[27];
assign P[17][28] = x[17] & y[28];
assign P[17][29] = x[17] & y[29];
assign P[17][30] = x[17] & y[30];
assign P[17][31] = x[17] & y[31];
assign P[18][0] = x[18] & y[0];
assign P[18][1] = x[18] & y[1];
assign P[18][2] = x[18] & y[2];
assign P[18][3] = x[18] & y[3];
assign P[18][4] = x[18] & y[4];
assign P[18][5] = x[18] & y[5];
assign P[18][6] = x[18] & y[6];
assign P[18][7] = x[18] & y[7];
assign P[18][8] = x[18] & y[8];
assign P[18][9] = x[18] & y[9];
assign P[18][10] = x[18] & y[10];
assign P[18][11] = x[18] & y[11];
assign P[18][12] = x[18] & y[12];
assign P[18][13] = x[18] & y[13];
assign P[18][14] = x[18] & y[14];
assign P[18][15] = x[18] & y[15];
assign P[18][16] = x[18] & y[16];
assign P[18][17] = x[18] & y[17];
assign P[18][18] = x[18] & y[18];
assign P[18][19] = x[18] & y[19];
assign P[18][20] = x[18] & y[20];
assign P[18][21] = x[18] & y[21];
assign P[18][22] = x[18] & y[22];
assign P[18][23] = x[18] & y[23];
assign P[18][24] = x[18] & y[24];
assign P[18][25] = x[18] & y[25];
assign P[18][26] = x[18] & y[26];
assign P[18][27] = x[18] & y[27];
assign P[18][28] = x[18] & y[28];
assign P[18][29] = x[18] & y[29];
assign P[18][30] = x[18] & y[30];
assign P[18][31] = x[18] & y[31];
assign P[19][0] = x[19] & y[0];
assign P[19][1] = x[19] & y[1];
assign P[19][2] = x[19] & y[2];
assign P[19][3] = x[19] & y[3];
assign P[19][4] = x[19] & y[4];
assign P[19][5] = x[19] & y[5];
assign P[19][6] = x[19] & y[6];
assign P[19][7] = x[19] & y[7];
assign P[19][8] = x[19] & y[8];
assign P[19][9] = x[19] & y[9];
assign P[19][10] = x[19] & y[10];
assign P[19][11] = x[19] & y[11];
assign P[19][12] = x[19] & y[12];
assign P[19][13] = x[19] & y[13];
assign P[19][14] = x[19] & y[14];
assign P[19][15] = x[19] & y[15];
assign P[19][16] = x[19] & y[16];
assign P[19][17] = x[19] & y[17];
assign P[19][18] = x[19] & y[18];
assign P[19][19] = x[19] & y[19];
assign P[19][20] = x[19] & y[20];
assign P[19][21] = x[19] & y[21];
assign P[19][22] = x[19] & y[22];
assign P[19][23] = x[19] & y[23];
assign P[19][24] = x[19] & y[24];
assign P[19][25] = x[19] & y[25];
assign P[19][26] = x[19] & y[26];
assign P[19][27] = x[19] & y[27];
assign P[19][28] = x[19] & y[28];
assign P[19][29] = x[19] & y[29];
assign P[19][30] = x[19] & y[30];
assign P[19][31] = x[19] & y[31];
assign P[20][0] = x[20] & y[0];
assign P[20][1] = x[20] & y[1];
assign P[20][2] = x[20] & y[2];
assign P[20][3] = x[20] & y[3];
assign P[20][4] = x[20] & y[4];
assign P[20][5] = x[20] & y[5];
assign P[20][6] = x[20] & y[6];
assign P[20][7] = x[20] & y[7];
assign P[20][8] = x[20] & y[8];
assign P[20][9] = x[20] & y[9];
assign P[20][10] = x[20] & y[10];
assign P[20][11] = x[20] & y[11];
assign P[20][12] = x[20] & y[12];
assign P[20][13] = x[20] & y[13];
assign P[20][14] = x[20] & y[14];
assign P[20][15] = x[20] & y[15];
assign P[20][16] = x[20] & y[16];
assign P[20][17] = x[20] & y[17];
assign P[20][18] = x[20] & y[18];
assign P[20][19] = x[20] & y[19];
assign P[20][20] = x[20] & y[20];
assign P[20][21] = x[20] & y[21];
assign P[20][22] = x[20] & y[22];
assign P[20][23] = x[20] & y[23];
assign P[20][24] = x[20] & y[24];
assign P[20][25] = x[20] & y[25];
assign P[20][26] = x[20] & y[26];
assign P[20][27] = x[20] & y[27];
assign P[20][28] = x[20] & y[28];
assign P[20][29] = x[20] & y[29];
assign P[20][30] = x[20] & y[30];
assign P[20][31] = x[20] & y[31];
assign P[21][0] = x[21] & y[0];
assign P[21][1] = x[21] & y[1];
assign P[21][2] = x[21] & y[2];
assign P[21][3] = x[21] & y[3];
assign P[21][4] = x[21] & y[4];
assign P[21][5] = x[21] & y[5];
assign P[21][6] = x[21] & y[6];
assign P[21][7] = x[21] & y[7];
assign P[21][8] = x[21] & y[8];
assign P[21][9] = x[21] & y[9];
assign P[21][10] = x[21] & y[10];
assign P[21][11] = x[21] & y[11];
assign P[21][12] = x[21] & y[12];
assign P[21][13] = x[21] & y[13];
assign P[21][14] = x[21] & y[14];
assign P[21][15] = x[21] & y[15];
assign P[21][16] = x[21] & y[16];
assign P[21][17] = x[21] & y[17];
assign P[21][18] = x[21] & y[18];
assign P[21][19] = x[21] & y[19];
assign P[21][20] = x[21] & y[20];
assign P[21][21] = x[21] & y[21];
assign P[21][22] = x[21] & y[22];
assign P[21][23] = x[21] & y[23];
assign P[21][24] = x[21] & y[24];
assign P[21][25] = x[21] & y[25];
assign P[21][26] = x[21] & y[26];
assign P[21][27] = x[21] & y[27];
assign P[21][28] = x[21] & y[28];
assign P[21][29] = x[21] & y[29];
assign P[21][30] = x[21] & y[30];
assign P[21][31] = x[21] & y[31];
assign P[22][0] = x[22] & y[0];
assign P[22][1] = x[22] & y[1];
assign P[22][2] = x[22] & y[2];
assign P[22][3] = x[22] & y[3];
assign P[22][4] = x[22] & y[4];
assign P[22][5] = x[22] & y[5];
assign P[22][6] = x[22] & y[6];
assign P[22][7] = x[22] & y[7];
assign P[22][8] = x[22] & y[8];
assign P[22][9] = x[22] & y[9];
assign P[22][10] = x[22] & y[10];
assign P[22][11] = x[22] & y[11];
assign P[22][12] = x[22] & y[12];
assign P[22][13] = x[22] & y[13];
assign P[22][14] = x[22] & y[14];
assign P[22][15] = x[22] & y[15];
assign P[22][16] = x[22] & y[16];
assign P[22][17] = x[22] & y[17];
assign P[22][18] = x[22] & y[18];
assign P[22][19] = x[22] & y[19];
assign P[22][20] = x[22] & y[20];
assign P[22][21] = x[22] & y[21];
assign P[22][22] = x[22] & y[22];
assign P[22][23] = x[22] & y[23];
assign P[22][24] = x[22] & y[24];
assign P[22][25] = x[22] & y[25];
assign P[22][26] = x[22] & y[26];
assign P[22][27] = x[22] & y[27];
assign P[22][28] = x[22] & y[28];
assign P[22][29] = x[22] & y[29];
assign P[22][30] = x[22] & y[30];
assign P[22][31] = x[22] & y[31];
assign P[23][0] = x[23] & y[0];
assign P[23][1] = x[23] & y[1];
assign P[23][2] = x[23] & y[2];
assign P[23][3] = x[23] & y[3];
assign P[23][4] = x[23] & y[4];
assign P[23][5] = x[23] & y[5];
assign P[23][6] = x[23] & y[6];
assign P[23][7] = x[23] & y[7];
assign P[23][8] = x[23] & y[8];
assign P[23][9] = x[23] & y[9];
assign P[23][10] = x[23] & y[10];
assign P[23][11] = x[23] & y[11];
assign P[23][12] = x[23] & y[12];
assign P[23][13] = x[23] & y[13];
assign P[23][14] = x[23] & y[14];
assign P[23][15] = x[23] & y[15];
assign P[23][16] = x[23] & y[16];
assign P[23][17] = x[23] & y[17];
assign P[23][18] = x[23] & y[18];
assign P[23][19] = x[23] & y[19];
assign P[23][20] = x[23] & y[20];
assign P[23][21] = x[23] & y[21];
assign P[23][22] = x[23] & y[22];
assign P[23][23] = x[23] & y[23];
assign P[23][24] = x[23] & y[24];
assign P[23][25] = x[23] & y[25];
assign P[23][26] = x[23] & y[26];
assign P[23][27] = x[23] & y[27];
assign P[23][28] = x[23] & y[28];
assign P[23][29] = x[23] & y[29];
assign P[23][30] = x[23] & y[30];
assign P[23][31] = x[23] & y[31];
assign P[24][0] = x[24] & y[0];
assign P[24][1] = x[24] & y[1];
assign P[24][2] = x[24] & y[2];
assign P[24][3] = x[24] & y[3];
assign P[24][4] = x[24] & y[4];
assign P[24][5] = x[24] & y[5];
assign P[24][6] = x[24] & y[6];
assign P[24][7] = x[24] & y[7];
assign P[24][8] = x[24] & y[8];
assign P[24][9] = x[24] & y[9];
assign P[24][10] = x[24] & y[10];
assign P[24][11] = x[24] & y[11];
assign P[24][12] = x[24] & y[12];
assign P[24][13] = x[24] & y[13];
assign P[24][14] = x[24] & y[14];
assign P[24][15] = x[24] & y[15];
assign P[24][16] = x[24] & y[16];
assign P[24][17] = x[24] & y[17];
assign P[24][18] = x[24] & y[18];
assign P[24][19] = x[24] & y[19];
assign P[24][20] = x[24] & y[20];
assign P[24][21] = x[24] & y[21];
assign P[24][22] = x[24] & y[22];
assign P[24][23] = x[24] & y[23];
assign P[24][24] = x[24] & y[24];
assign P[24][25] = x[24] & y[25];
assign P[24][26] = x[24] & y[26];
assign P[24][27] = x[24] & y[27];
assign P[24][28] = x[24] & y[28];
assign P[24][29] = x[24] & y[29];
assign P[24][30] = x[24] & y[30];
assign P[24][31] = x[24] & y[31];
assign P[25][0] = x[25] & y[0];
assign P[25][1] = x[25] & y[1];
assign P[25][2] = x[25] & y[2];
assign P[25][3] = x[25] & y[3];
assign P[25][4] = x[25] & y[4];
assign P[25][5] = x[25] & y[5];
assign P[25][6] = x[25] & y[6];
assign P[25][7] = x[25] & y[7];
assign P[25][8] = x[25] & y[8];
assign P[25][9] = x[25] & y[9];
assign P[25][10] = x[25] & y[10];
assign P[25][11] = x[25] & y[11];
assign P[25][12] = x[25] & y[12];
assign P[25][13] = x[25] & y[13];
assign P[25][14] = x[25] & y[14];
assign P[25][15] = x[25] & y[15];
assign P[25][16] = x[25] & y[16];
assign P[25][17] = x[25] & y[17];
assign P[25][18] = x[25] & y[18];
assign P[25][19] = x[25] & y[19];
assign P[25][20] = x[25] & y[20];
assign P[25][21] = x[25] & y[21];
assign P[25][22] = x[25] & y[22];
assign P[25][23] = x[25] & y[23];
assign P[25][24] = x[25] & y[24];
assign P[25][25] = x[25] & y[25];
assign P[25][26] = x[25] & y[26];
assign P[25][27] = x[25] & y[27];
assign P[25][28] = x[25] & y[28];
assign P[25][29] = x[25] & y[29];
assign P[25][30] = x[25] & y[30];
assign P[25][31] = x[25] & y[31];
assign P[26][0] = x[26] & y[0];
assign P[26][1] = x[26] & y[1];
assign P[26][2] = x[26] & y[2];
assign P[26][3] = x[26] & y[3];
assign P[26][4] = x[26] & y[4];
assign P[26][5] = x[26] & y[5];
assign P[26][6] = x[26] & y[6];
assign P[26][7] = x[26] & y[7];
assign P[26][8] = x[26] & y[8];
assign P[26][9] = x[26] & y[9];
assign P[26][10] = x[26] & y[10];
assign P[26][11] = x[26] & y[11];
assign P[26][12] = x[26] & y[12];
assign P[26][13] = x[26] & y[13];
assign P[26][14] = x[26] & y[14];
assign P[26][15] = x[26] & y[15];
assign P[26][16] = x[26] & y[16];
assign P[26][17] = x[26] & y[17];
assign P[26][18] = x[26] & y[18];
assign P[26][19] = x[26] & y[19];
assign P[26][20] = x[26] & y[20];
assign P[26][21] = x[26] & y[21];
assign P[26][22] = x[26] & y[22];
assign P[26][23] = x[26] & y[23];
assign P[26][24] = x[26] & y[24];
assign P[26][25] = x[26] & y[25];
assign P[26][26] = x[26] & y[26];
assign P[26][27] = x[26] & y[27];
assign P[26][28] = x[26] & y[28];
assign P[26][29] = x[26] & y[29];
assign P[26][30] = x[26] & y[30];
assign P[26][31] = x[26] & y[31];
assign P[27][0] = x[27] & y[0];
assign P[27][1] = x[27] & y[1];
assign P[27][2] = x[27] & y[2];
assign P[27][3] = x[27] & y[3];
assign P[27][4] = x[27] & y[4];
assign P[27][5] = x[27] & y[5];
assign P[27][6] = x[27] & y[6];
assign P[27][7] = x[27] & y[7];
assign P[27][8] = x[27] & y[8];
assign P[27][9] = x[27] & y[9];
assign P[27][10] = x[27] & y[10];
assign P[27][11] = x[27] & y[11];
assign P[27][12] = x[27] & y[12];
assign P[27][13] = x[27] & y[13];
assign P[27][14] = x[27] & y[14];
assign P[27][15] = x[27] & y[15];
assign P[27][16] = x[27] & y[16];
assign P[27][17] = x[27] & y[17];
assign P[27][18] = x[27] & y[18];
assign P[27][19] = x[27] & y[19];
assign P[27][20] = x[27] & y[20];
assign P[27][21] = x[27] & y[21];
assign P[27][22] = x[27] & y[22];
assign P[27][23] = x[27] & y[23];
assign P[27][24] = x[27] & y[24];
assign P[27][25] = x[27] & y[25];
assign P[27][26] = x[27] & y[26];
assign P[27][27] = x[27] & y[27];
assign P[27][28] = x[27] & y[28];
assign P[27][29] = x[27] & y[29];
assign P[27][30] = x[27] & y[30];
assign P[27][31] = x[27] & y[31];
assign P[28][0] = x[28] & y[0];
assign P[28][1] = x[28] & y[1];
assign P[28][2] = x[28] & y[2];
assign P[28][3] = x[28] & y[3];
assign P[28][4] = x[28] & y[4];
assign P[28][5] = x[28] & y[5];
assign P[28][6] = x[28] & y[6];
assign P[28][7] = x[28] & y[7];
assign P[28][8] = x[28] & y[8];
assign P[28][9] = x[28] & y[9];
assign P[28][10] = x[28] & y[10];
assign P[28][11] = x[28] & y[11];
assign P[28][12] = x[28] & y[12];
assign P[28][13] = x[28] & y[13];
assign P[28][14] = x[28] & y[14];
assign P[28][15] = x[28] & y[15];
assign P[28][16] = x[28] & y[16];
assign P[28][17] = x[28] & y[17];
assign P[28][18] = x[28] & y[18];
assign P[28][19] = x[28] & y[19];
assign P[28][20] = x[28] & y[20];
assign P[28][21] = x[28] & y[21];
assign P[28][22] = x[28] & y[22];
assign P[28][23] = x[28] & y[23];
assign P[28][24] = x[28] & y[24];
assign P[28][25] = x[28] & y[25];
assign P[28][26] = x[28] & y[26];
assign P[28][27] = x[28] & y[27];
assign P[28][28] = x[28] & y[28];
assign P[28][29] = x[28] & y[29];
assign P[28][30] = x[28] & y[30];
assign P[28][31] = x[28] & y[31];
assign P[29][0] = x[29] & y[0];
assign P[29][1] = x[29] & y[1];
assign P[29][2] = x[29] & y[2];
assign P[29][3] = x[29] & y[3];
assign P[29][4] = x[29] & y[4];
assign P[29][5] = x[29] & y[5];
assign P[29][6] = x[29] & y[6];
assign P[29][7] = x[29] & y[7];
assign P[29][8] = x[29] & y[8];
assign P[29][9] = x[29] & y[9];
assign P[29][10] = x[29] & y[10];
assign P[29][11] = x[29] & y[11];
assign P[30][31] = x[30] & y[31];
assign P[31][0] = x[31] & y[0];
assign P[31][1] = x[31] & y[1];
assign P[31][2] = x[31] & y[2];
assign P[31][3] = x[31] & y[3];
assign P[31][4] = x[31] & y[4];
assign P[31][5] = x[31] & y[5];
assign P[31][6] = x[31] & y[6];
assign P[31][7] = x[31] & y[7];
assign P[31][8] = x[31] & y[8];
assign P[31][9] = x[31] & y[9];
assign P[31][10] = x[31] & y[10];
assign P[31][11] = x[31] & y[11];
assign P[31][12] = x[31] & y[12];
assign P[31][13] = x[31] & y[13];
assign P[31][14] = x[31] & y[14];
assign P[31][15] = x[31] & y[15];
assign P[31][16] = x[31] & y[16];
assign P[31][17] = x[31] & y[17];
assign P[31][18] = x[31] & y[18];
assign P[31][19] = x[31] & y[19];
assign P[31][20] = x[31] & y[20];
assign P[31][21] = x[31] & y[21];
assign P[31][22] = x[31] & y[22];
assign P[31][23] = x[31] & y[23];
assign P[31][24] = x[31] & y[24];
assign P[31][25] = x[31] & y[25];
assign P[31][26] = x[31] & y[26];
assign P[31][27] = x[31] & y[27];
assign P[31][28] = x[31] & y[28];
assign P[31][29] = x[31] & y[29];
assign P[31][30] = x[31] & y[30];
assign P[31][31] = x[31] & y[31];


assign P[29][12] = x[29] & y[12];
assign P[29][13] = x[29] & y[13];
assign P[29][14] = x[29] & y[14];
assign P[29][15] = x[29] & y[15];
assign P[29][16] = x[29] & y[16];
assign P[29][17] = x[29] & y[17];
assign P[29][18] = x[29] & y[18];
assign P[29][19] = x[29] & y[19];
assign P[29][20] = x[29] & y[20];
assign P[29][21] = x[29] & y[21];
assign P[29][22] = x[29] & y[22];
assign P[29][23] = x[29] & y[23];
assign P[29][24] = x[29] & y[24];
assign P[29][25] = x[29] & y[25];
assign P[29][26] = x[29] & y[26];
assign P[29][27] = x[29] & y[27];
assign P[29][28] = x[29] & y[28];
assign P[29][29] = x[29] & y[29];
assign P[29][30] = x[29] & y[30];
assign P[29][31] = x[29] & y[31];
assign P[30][0] = x[30] & y[0];
assign P[30][1] = x[30] & y[1];
assign P[30][2] = x[30] & y[2];
assign P[30][3] = x[30] & y[3];
assign P[30][4] = x[30] & y[4];
assign P[30][5] = x[30] & y[5];
assign P[30][6] = x[30] & y[6];
assign P[30][7] = x[30] & y[7];
assign P[30][8] = x[30] & y[8];
assign P[30][9] = x[30] & y[9];
assign P[30][10] = x[30] & y[10];
assign P[30][11] = x[30] & y[11];
assign P[30][12] = x[30] & y[12];
assign P[30][13] = x[30] & y[13];
assign P[30][14] = x[30] & y[14];
assign P[30][15] = x[30] & y[15];
assign P[30][16] = x[30] & y[16];
assign P[30][17] = x[30] & y[17];
assign P[30][18] = x[30] & y[18];
assign P[30][19] = x[30] & y[19];
assign P[30][20] = x[30] & y[20];
assign P[30][21] = x[30] & y[21];
assign P[30][22] = x[30] & y[22];
assign P[30][23] = x[30] & y[23];
assign P[30][24] = x[30] & y[24];
assign P[30][25] = x[30] & y[25];
assign P[30][26] = x[30] & y[26];
assign P[30][27] = x[30] & y[27];
assign P[30][28] = x[30] & y[28];
assign P[30][29] = x[30] & y[29];
assign P[30][30] = x[30] & y[30];
assign P[30][31] = x[30] & y[31];
assign P[31][0] = x[31] & y[0];
assign P[31][1] = x[31] & y[1];
assign P[31][2] = x[31] & y[2];
assign P[31][3] = x[31] & y[3];
assign P[31][4] = x[31] & y[4];
assign P[31][5] = x[31] & y[5];
assign P[31][6] = x[31] & y[6];
assign P[31][7] = x[31] & y[7];
assign P[31][8] = x[31] & y[8];
assign P[31][9] = x[31] & y[9];
assign P[31][10] = x[31] & y[10];
assign P[31][11] = x[31] & y[11];
assign P[31][12] = x[31] & y[12];
assign P[31][13] = x[31] & y[13];
assign P[31][14] = x[31] & y[14];
assign P[31][15] = x[31] & y[15];
assign P[31][16] = x[31] & y[16];
assign P[31][17] = x[31] & y[17];
assign P[31][18] = x[31] & y[18];
assign P[31][19] = x[31] & y[19];
assign P[31][20] = x[31] & y[20];
assign P[31][21] = x[31] & y[21];
assign P[31][22] = x[31] & y[22];
assign P[31][23] = x[31] & y[23];
assign P[31][24] = x[31] & y[24];
assign P[31][25] = x[31] & y[25];
assign P[31][26] = x[31] & y[26];
assign P[31][27] = x[31] & y[27];
assign P[31][28] = x[31] & y[28];
assign P[31][29] = x[31] & y[29];
assign P[31][30] = x[31] & y[30];
assign P[31][31] = x[31] & y[31];

wire [63:0] s[63:0];
genvar p1;
for(p1=0;p1<32;p1=p1+1)begin
assign s[0][p1]=P[0][p1];
assign s[1][p1+1]=P[1][p1];
assign s[2][p1+2]=P[2][p1];
assign s[3][p1+3]=P[3][p1];
assign s[4][p1+4]=P[4][p1];
assign s[5][p1+5]=P[5][p1];
assign s[6][p1+6]=P[6][p1];
assign s[7][p1+7]=P[7][p1];
assign s[8][p1+8]=P[8][p1];
assign s[9][p1+9]=P[9][p1];
assign s[10][p1+10]=P[10][p1];
assign s[11][p1+11]=P[11][p1];
assign s[12][p1+12]=P[12][p1];
assign s[13][p1+13]=P[13][p1];
assign s[14][p1+14]=P[14][p1];
assign s[15][p1+15]=P[15][p1];
assign s[16][p1+16]=P[16][p1];
assign s[17][p1+17]=P[17][p1];
assign s[18][p1+18]=P[18][p1];
assign s[19][p1+19]=P[19][p1];
assign s[20][p1+20]=P[20][p1];
assign s[21][p1+21]=P[21][p1];
assign s[22][p1+22]=P[22][p1];
assign s[23][p1+23]=P[23][p1];
assign s[24][p1+24]=P[24][p1];
assign s[25][p1+25]=P[25][p1];
assign s[26][p1+26]=P[26][p1];
assign s[27][p1+27]=P[27][p1];
assign s[28][p1+28]=P[28][p1];
assign s[29][p1+29]=P[29][p1];
assign s[30][p1+30]=P[30][p1];
assign s[31][p1+31]=P[31][p1];
end

genvar p2;
for(p2=32;p2<64;p2=p2+1)begin
assign s[0][p2]=1'b0;
assign s[1][p2+1]=1'b0;
assign s[2][p2+2]=1'b0;
assign s[3][p2+3]=1'b0;
assign s[4][p2+4]=1'b0;
assign s[5][p2+5]=1'b0;
assign s[6][p2+6]=1'b0;
assign s[7][p2+7]=1'b0;
assign s[8][p2+8]=1'b0;
assign s[9][p2+9]=1'b0;
assign s[10][p2+10]=1'b0;
assign s[11][p2+11]=1'b0;
assign s[12][p2+12]=1'b0;
assign s[13][p2+13]=1'b0;
assign s[14][p2+14]=1'b0;
assign s[15][p2+15]=1'b0;
assign s[16][p2+16]=1'b0;
assign s[17][p2+17]=1'b0;
assign s[18][p2+18]=1'b0;
assign s[19][p2+19]=1'b0;
assign s[20][p2+20]=1'b0;
assign s[21][p2+21]=1'b0;
assign s[22][p2+22]=1'b0;
assign s[23][p2+23]=1'b0;
assign s[24][p2+24]=1'b0;
assign s[25][p2+25]=1'b0;
assign s[26][p2+26]=1'b0;
assign s[27][p2+27]=1'b0;
assign s[28][p2+28]=1'b0;
assign s[29][p2+29]=1'b0;
assign s[30][p2+30]=1'b0;
assign s[31][p2+31]=1'b0;
end
genvar p3;



assign s[1][0]=1'b0;
assign s[2][1:0]=2'b00;
assign s[3][2:0]=3'b000;
assign s[4][3:0]=4'b0000;
assign s[5][4:0]=5'b00000;
assign s[6][5:0]=6'b000000;
assign s[7][6:0]=7'b0000000;
assign s[8][7:0]=8'b00000000;
assign s[9][8:0]=9'b000000000;
assign s[10][9:0]=10'b0000000000;
assign s[11][10:0]=11'b00000000000;
assign s[12][11:0]=12'b000000000000;
assign s[13][12:0]=13'b0000000000000;
assign s[14][13:0]=14'b00000000000000;
assign s[15][14:0]=15'b000000000000000;
assign s[16][15:0]=16'b0000000000000000;
assign s[17][16:0]=17'b00000000000000000;
assign s[18][17:0]=18'b000000000000000000;
assign s[19][18:0]=19'b0000000000000000000;
assign s[20][19:0]=20'b00000000000000000000;
assign s[21][20:0]=21'b000000000000000000000;
assign s[22][21:0]=22'b0000000000000000000000;
assign s[23][22:0]=23'b00000000000000000000000;
assign s[24][23:0]=24'b000000000000000000000000;
assign s[25][24:0]=25'b0000000000000000000000000;
assign s[26][25:0]=26'b00000000000000000000000000;
assign s[27][26:0]=27'b000000000000000000000000000;
assign s[28][27:0]=28'b0000000000000000000000000000;
assign s[29][28:0]=29'b00000000000000000000000000000;
assign s[30][29:0]=30'b000000000000000000000000000000;
assign s[31][30:0]=31'b0000000000000000000000000000000;


wire [63:0]s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,cout;

adder64bit u1 (s[0][63:0],s[1][63:0],s1[63:0]);
adder64bit u2 (s[2][63:0],s1,s2);
adder64bit u3 (s[3][63:0],s2,s3);
adder64bit u4 (s[4][63:0],s3,s4);
adder64bit u5 (s[5][63:0],s4,s5);
adder64bit u6 (s[6][63:0],s5,s6);
adder64bit u7 (s[7][63:0],s6,s7);
adder64bit u8 (s[8][63:0],s7,s8);
adder64bit u9 (s[9][63:0],s8,s9);
adder64bit u10 (s[10][63:0],s9,s10);
adder64bit u11 (s[11][63:0],s10,s11);
adder64bit u12 (s[12][63:0],s11,s12);
adder64bit u13(s[13][63:0],s12,s13);
adder64bit u14 (s [14][63:0],s13,s14);
adder64bit u15(s[15][63:0],s14,s15);
adder64bit u16(s[16][63:0],s15,s16);
adder64bit u17 (s[17][63:0],s16,s17);
adder64bit u18 (s[18][63:0],s17,s18);
adder64bit  u19 (s[19][63:0],s18,s19);
adder64bit u20 (s[20][63:0],s19,s20);
adder64bit u21(s[21][63:0],s20,s21);
adder64bit u22 (s[22][63:0],s21,s22);
adder64bit u23 (s[23][63:0],s22,s23);
adder64bit u24( s[24][63:0],s23,s24);
adder64bit u25 (s[25][63:0],s24,s25);
adder64bit u26 (s[26][63:0],s25,s26);
adder64bit u27 (s[27][63:0],s26,s27);
adder64bit u28 (s[28][63:0],s27,s28);
adder64bit u29 (s[29][63:0],s28,s29);
adder64bit u30 (s[30][63:0],s29,s30);
adder64bit u31 (s[31][63:0],s30,cout);

assign z = cout;


endmodule

